LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;

ENTITY FFD IS
	PORT(
		D, CLK, RST:IN STD_LOGIC;
		Q: OUT STD_LOGIC);
END FFD;

ARCHITECTURE arch OF FFD IS
BEGIN
	PROCESS(CLK)
	BEGIN
		IF RST='0' THEN 
				Q <= '0';
		ELSIF RISING_EDGE(CLK) THEN 
				Q <= D;
		END IF;
		
	END PROCESS;
END arch;